module elevator